// File: alucodes.sv
// Author: Tommy Sætre
// Description: Constants defining alu codes for readability in alu source code
// Last revision: 27/02/24
// **AI NOTICE: Directly copied from code written by T. Kazmierski.

`define RA      3'b000
`define RB      3'b001
`define RADD    3'b010
`define RSUB    3'b011
`define RAND    3'b100
`define ROR     3'b101
`define RXOR    3'b110
`define RMUL    3'b111